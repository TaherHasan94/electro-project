* C:\Users\User\Desktop\Project Electro\Thermistor\Yazan&Taher&AhmadProject.sch

* Schematics Version 9.1 - Web Update 1
* Fri Jun 17 16:07:55 2022


.PARAM         Rs=40k 

** Analysis setup **
.DC LIN PARAM Rs 40k 10k 500 
.tran 0ns 1000ns
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Yazan&Taher&AhmadProject.net"
.INC "Yazan&Taher&AhmadProject.als"


.probe


.END
